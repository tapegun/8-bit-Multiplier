module Processor()