module register_unit()